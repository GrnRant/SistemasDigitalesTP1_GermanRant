library IEEE;
use IEEE.std_logic_1164.all;

package semaforos_states is
    type semf_states is (E0, E1, E2, E3, E4 , E5);
end package semaforos_states;
